*Cmos Inverter involving equating Rise and Fall Time
**Including suitable model definition files
.include model.txt 
**Variables to be used in program
.param lambda=90n	
.param Wn=0.6u
.param Wp=1.55795u 

**name D G S B type length width  area of source  perimeter of source  area of drain   perimeter of drain-------------------- 
***------------------------------------- NMOS-----------------------------------------------------------------------------***


m_n1 o1 input 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n2 in_DUT o1 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_DUT in_Fan in_DUT 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout1 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout2 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout3 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout4 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout5 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout6 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout7 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}
m_n_Fanout8 output in_Fan 0 0 cmosn L=0.4u W=Wn AS={4*lambda*Wn} PS={2*Wn+8*lambda} AD={4*lambda*Wn} PD={2*Wn+8*lambda}

****-------------------------------------PMOS----------------------------------------------------------------------------****
m_p1 o1 input sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p2 in_DUT o1 sup sup cmosp L=0.4u  W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_DUT in_Fan in_DUT sup sup cmosp L=0.4u  W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout1 output in_Fan sup sup cmosp L=0.4u  W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout2 output in_Fan sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout3 output in_Fan sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout4 output in_Fan sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout5 output in_Fan sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout6 output in_Fan sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout7 output in_Fan sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}
m_p_Fanout8 output in_Fan sup sup cmosp L=0.4u W=Wp AS={4*lambda*Wp} PS={2*Wp+8*lambda} AD={4*lambda*Wp} PD={2*Wp+8*lambda}



**Attaching the load.........................................................................................................
C_load output 0 0.1p
	
**Defining Supply............................................................................................................
Vdd sup 0 dc 3.3v	

**Setting Up the input pulse –----------------------------------------------------------------------------------------------
** pulse(<initial value> <pulsed value> <Timedelay> <risetime> <falltime> <pulsewidth> <period>)**
vin input 0 pulse(0 3.3 0 0.5p 0.5p 0.1u 0.2u)

**Running Transient analysis –-----------------------------------------------------------------------------------------------
*** .tran <tstep> <tstop> ***
.tran 1p 1us

**Measurement of rise time and fall time –-----------------------------------------------------------------------------------

*.measure tran rise_output trig v(output) val=0.33 rise=1 targ v(output) val=2.97 rise=1
*.measure tran fall_output trig v(output) val=2.97 fall=1 targ v(output) val=0.33 fall=1

*.measure tran rise_DUT trig v(in_Fan) val=0.33 rise=1 targ v(in_Fan) val=2.97 rise=1
*.measure tran fall_DUT trig v(in_Fan) val=2.97 fall=1 targ v(in_Fan) val=0.33 fall=1
.measure tran delay_DUT trig v(in_DUT) val=1.65 rise=1 targ v(in_Fan) val=1.65 fall=1

**Output plotting –----------------------------------------------------------------------------------------------------------
.control
run
plot v(in_DUT) v(in_Fan)
**hardcopy [file name] [plot arguments]
**gnuplot delay v(in_DUT) v(in_Fan) 
**gnuplot inout v(input) v(output)
.endc
.end

